module Comb_Assign (
    input wire in2,
    output wire out,
    input wire in1
);
    assign out = in1 & in2;
endmodule

