module coalesced_assign (
    input logic [3:0] in_l,
    output logic [7:0] out,
    input logic [3:0] in_h
);
    wire [7:0] temp_wire;
    assign temp_wire[7:4] = in_h;
    assign temp_wire[3:0] = in_l;
    assign out = temp_wire;
endmodule

