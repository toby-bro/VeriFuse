module multi_always_comb (
    output wire [7:0] out1,
    output wire [7:0] out2,
    input wire [7:0] in1,
    input wire [7:0] in2
);
    logic [7:0] intermediate1;
    logic [7:0] intermediate2;
    always @(*) begin
        intermediate1 = in1 & in2;
    end
    always @(*) begin
        intermediate2 = in1 | in2;
    end
    assign out1 = intermediate1 + 8'd1;
    assign out2 = intermediate2 - 8'd1;
endmodule

