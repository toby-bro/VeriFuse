module simple_logic_b (
    output wire data_d,
    input wire data_c
);
    assign data_d = data_c;
endmodule

