module SequentialLogicPlaceholder (
    input logic clk,
    input logic rst,
    input logic [15:0] data_in,
    output logic [15:0] data_out
);
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            data_out <= 16'h0;
        end else begin
            data_out <= data_in;
        end
    end
endmodule

