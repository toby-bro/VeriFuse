module split_input_only_var (
    input logic [7:0] data_in_k,
    output logic [7:0] data_out_k,
    input logic clk_k,
    input logic control_signal_k
);
    always @(posedge clk_k) begin
       if (control_signal_k) begin
          data_out_k <= data_in_k;
       end
    end
endmodule

