interface my_if;
    logic valid;
    logic [7:0] data;
    logic ready;

    modport FullAccess (
        input data,
        input output ready,
        input output valid
    );

    modport AccessIn (
        output data,
        output output valid,
        output input ready
    );

    modport AccessOut (
        input data,
        input input valid,
        input output ready
    );

    logic [7:0] data;
      logic ready;
      logic valid;
      modport FullAccess (input data, output ready, output valid);
      modport AccessIn (output data, output valid, input ready);
      modport AccessOut (input data, input valid, output ready);
endinterface
module module_case_write (
    input logic [1:0] select_case,
    input logic [7:0] data_case_a,
    input logic [7:0] data_case_b,
    output logic case_output_ready
);
    my_if case_vif_inst();
      always_comb begin
    case (select_case)
      2'b00: begin
        case_vif_inst.data = 8'hAA;
        case_vif_inst.valid = 1'b1;
        case_vif_inst.ready = 1'b0;
      end
      2'b01: begin
        case_vif_inst.data = data_case_a;
        case_vif_inst.valid = 1'b0;
        case_vif_inst.ready = 1'b1;
      end
      2'b10: begin
        case_vif_inst.data = data_case_b;
        case_vif_inst.valid = 1'b1;
        case_vif_inst.ready = 1'b1;
      end
      default: begin
        case_vif_inst.data = 8'hFF;
        case_vif_inst.valid = 1'b0;
        case_vif_inst.ready = 1'b0;
      end
    endcase
    case_output_ready = case_vif_inst.ready;
      end
endmodule

