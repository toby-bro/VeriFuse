module dup_literal_param (
    output logic [7:0] final_result,
    input logic [4:0] index
);
    parameter CONST_A = 8'd10;
    localparam CONST_B = 8'd20;
    parameter CONST_C = 10;
    localparam CONST_D = 8'hFF;
    parameter CONST_E = 8'b01010101;
    logic [7:0] temp1, temp2;
    assign temp1 = index + CONST_A;
    assign temp2 = index + 10;
    always_comb begin
        logic [7:0] local_temp;
        local_temp = index * CONST_B;
        final_result = temp1 + temp2 + local_temp;
        if (index > 5) begin
            final_result = final_result + 1;
        end else if (index < CONST_C) begin
            final_result = final_result - 1;
        end
        case (index)
            5'd0: final_result = CONST_A;
            5'd1: final_result = 20;
            5'd2: final_result = 10;
            5'd3: final_result = CONST_B;
            5'd4: final_result = CONST_D;
            5'd5: final_result = 8'hFF;
            default: final_result = CONST_E;
        endcase
    end
endmodule

