interface my_if;
    logic valid;
    logic [7:0] data;
    logic ready;

    modport FullAccess (
        input data,
        input output ready,
        input output valid
    );

    modport AccessIn (
        output data,
        output output valid,
        output input ready
    );

    modport AccessOut (
        input data,
        input input valid,
        input output ready
    );

    logic [7:0] data;
      logic ready;
      logic valid;
      modport FullAccess (input data, output ready, output valid);
      modport AccessIn (output data, output valid, input ready);
      modport AccessOut (input data, input valid, output ready);
endinterface
module module_task_write (
    input logic task_en,
    input logic [7:0] in_task_data,
    output logic task_output_valid
);
    my_if task_vif_inst();
      task automatic update_vif_signals(input logic en, input logic [7:0] data_val,
                                    output logic [7:0] vif_data, output logic vif_valid, output logic vif_ready);
    if (en) begin
      vif_data = data_val;
      vif_valid = 1'b1;
      vif_ready = 1'b0;
    end else begin
      vif_data = 8'h0;
      vif_valid = 1'b0;
      vif_ready = 1'b1;
    end
      endtask
      always_comb begin
    update_vif_signals(task_en, in_task_data, task_vif_inst.data, task_vif_inst.valid, task_vif_inst.ready);
    task_output_valid = task_vif_inst.valid;
      end
endmodule

