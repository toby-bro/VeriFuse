module mismatched_width_unhandled (
    input logic [7:0] in,
    output logic [3:0] out
);
    assign out = in;
endmodule

