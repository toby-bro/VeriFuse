module more_procedural (
    input logic [31:0] p_in1,
    input logic [31:0] p_in2,
    output logic [31:0] p_out,
    input logic [1:0] p_mode
);
    always_comb begin
    case (p_mode)
      2'b00: p_out = (p_in1 + p_in2) * 2;
      2'b01: p_out = (p_in1 - p_in2) / 3; 
      2'b10: p_out = (p_in1 << 4) | (p_in2 >> 2);
      default: p_out = ~(p_in1 ^ p_in2) + 1;
    endcase
      end
endmodule

