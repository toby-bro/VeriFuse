module simple_and_gate (
    output logic out,
    input logic in1,
    input logic in2
);
    assign out = in1 & in2;
endmodule

