../testbench.sv