module keyword_import_export (
    input logic keyword_in,
    output logic keyword_out
);
    assign keyword_out = keyword_in;
endmodule

