module SimpleAssign (
    output logic [9:0] val_out,
    input logic [9:0] val_in
);
    assign val_out = val_in;
endmodule

