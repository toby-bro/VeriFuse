module loop_with_internal_assign (
    output logic [7:0] final_val,
    input logic [3:0] start_val
);
    logic [7:0] current_val;
      always_comb begin
    current_val = start_val;
    for (int k = 0; k < 3; k = k + 1) begin
      current_val = current_val + 1;
    end
    final_val = current_val;
      end
endmodule

