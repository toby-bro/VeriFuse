module split_vector_assign (
    input logic condition_y,
    input logic [7:0] in_val_y,
    output logic [7:0] out_vec_y,
    input logic clk_y
);
    always @(posedge clk_y) begin
        if (condition_y) begin
            out_vec_y[3:0] <= in_val_y[3:0];
            out_vec_y[7:4] <= in_val_y[7:4] + 1;
        end else begin
            out_vec_y <= 8'hFF;
        end
    end
endmodule

