module split_mixed_cond_seq (
    input logic condition_e,
    input logic [7:0] in_val_e,
    input logic [7:0] in_override_e,
    output logic [7:0] out_val_e,
    output logic status_e,
    input logic clk_e
);
    logic [7:0] temp_val_e;
    always @(posedge clk_e) begin
        temp_val_e <= in_val_e + 5;
        if (condition_e) begin
            out_val_e <= temp_val_e;
            status_e <= 1;
        end else begin
            out_val_e <= in_override_e;
            status_e <= 0;
        end
    end
endmodule

