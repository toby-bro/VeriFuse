module keyword_import_export (
    output logic keyword_out,
    input logic keyword_in
);
    assign keyword_out = keyword_in;
endmodule

