module ArrayIndexAndPartSelect (
    input logic [4:0] start_bit,
    output logic bit_out,
    output logic [7:0] byte_out,
    input logic [31:0] data_in,
    input int index_in
);
    logic [31:0] internal_data = data_in;
    assign bit_out = internal_data[index_in];
    assign byte_out = internal_data[start_bit +: 8];
endmodule

