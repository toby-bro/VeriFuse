/home/jns/Documents/Berkeley/ibex/rtl/ibex_branch_predict.sv