module simple_xor_gate (
    input logic in2,
    output logic out,
    input logic in1
);
    assign out = in1 ^ in2;
endmodule

